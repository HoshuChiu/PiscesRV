module ifu_decoder (
    input wire [31:0] ;
);

endmodule //ifu_decoder